module //name //(port list);
	//data type declarations
	//functionality statements
	//timing specifications

endmodule